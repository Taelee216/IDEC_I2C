module asbc();

endmodule