module asbc();
    asdasdf
    asdfasd
    asdfasdf
    
endmodule